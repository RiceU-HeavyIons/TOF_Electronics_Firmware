two_by_3bit_mux_inst : two_by_3bit_mux PORT MAP (
		data1x	 => data1x_sig,
		data0x	 => data0x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
