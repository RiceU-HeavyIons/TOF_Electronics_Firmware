bus_tri_8_inst : bus_tri_8 PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		enabletr	 => enabletr_sig,
		tridata	 => tridata_sig,
		result	 => result_sig
	);
