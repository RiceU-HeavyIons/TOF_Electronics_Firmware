mux_4_to_1_1bit_inst : mux_4_to_1_1bit PORT MAP (
		data3	 => data3_sig,
		data2	 => data2_sig,
		data1	 => data1_sig,
		data0	 => data0_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
