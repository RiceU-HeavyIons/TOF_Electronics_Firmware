TFF_LB_inst : TFF_LB PORT MAP (
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);
