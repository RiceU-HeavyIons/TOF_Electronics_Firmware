mux_2_to_1_3bit_inst : mux_2_to_1_3bit PORT MAP (
		data1x	 => data1x_sig,
		data0x	 => data0x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
