mux_2x32_inst : mux_2x32 PORT MAP (
		data1x	 => data1x_sig,
		data0x	 => data0x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
