ctr12bit_inst : ctr12bit PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
