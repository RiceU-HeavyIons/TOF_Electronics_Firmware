dff_sclr_sset_inst : dff_sclr_sset PORT MAP (
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		sset	 => sset_sig,
		data	 => data_sig,
		q	 => q_sig
	);
