-- $Id: serdes_reader.vhd,v 1.5 2007-12-27 20:23:15 jschamba Exp $
-------------------------------------------------------------------------------
-- Title      : Serdes Reader
-- Project    : 
-------------------------------------------------------------------------------
-- File       : serdes_reader.vhd
-- Author     : 
-- Company    : 
-- Created    : 2007-11-21
-- Last update: 2007-12-27
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Reads the data from the Serdes FPGA and generates the
--              necessary signals to latch it into a (dual clock) FIFO
-------------------------------------------------------------------------------
-- Copyright (c) 2007 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2007-11-21  1.0      jschamba        Created
-------------------------------------------------------------------------------


LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.ALL;
LIBRARY lpm;
USE lpm.lpm_components.ALL;
LIBRARY altera;
USE altera.altera_primitives_components.ALL;
USE work.my_conversions.ALL;
USE work.my_utilities.ALL;

ENTITY serdes_reader IS
  
  PORT (
    clk80mhz            : IN  std_logic;
    areset_n            : IN  std_logic;
    indata              : IN  std_logic_vector(15 DOWNTO 0);
    fifo_empty          : IN  std_logic;
    outfifo_almost_full : IN  boolean;
    evt_trg             : IN  std_logic;
    trgFifo_empty       : IN  std_logic;
    trgFifo_q           : IN  std_logic_vector (19 DOWNTO 0);
    trgFifo_rdreq       : OUT std_logic;
    busy                : OUT std_logic;  -- active low
    rdsel_out           : OUT std_logic_vector(1 DOWNTO 0);
    rdreq_out           : OUT std_logic;
    wrreq_out           : OUT std_logic;  -- assuming FIFO clk is clk80mhz
    outdata             : OUT std_logic_vector(31 DOWNTO 0)
    );

END ENTITY serdes_reader;

ARCHITECTURE a OF serdes_reader IS

  SIGNAL s_outdata   : std_logic_vector (31 DOWNTO 0);
  SIGNAL s_wrreq_out : std_logic;

  TYPE TState_type IS (
    SWaitTrig,
    SFifoChk,
    STagWrd,
    SRdSerA,
    SDelay,
    SRdTrg,
    SEnd
    );
  SIGNAL TState : TState_type;
  
BEGIN  -- ARCHITECTURE a

  rdsel_out <= "00";
  wrreq_out <= s_wrreq_out;
  outdata   <= s_outdata;


  shifter : PROCESS (clk80mhz, areset_n) IS
    VARIABLE ctr       : integer RANGE 0 TO 2    := 0;
    VARIABLE delayCtr  : integer RANGE 0 TO 2047 := 0;
    VARIABLE block_end : boolean;
  BEGIN
    IF areset_n = '0' THEN              -- asynchronous reset (active low)
      s_outdata     <= (OTHERS => '0');
      ctr           := 0;
      rdreq_out     <= '0';
      block_end     := false;
      TState        <= SWaitTrig;
      busy          <= '0';             -- default is "busy"
      trgFifo_rdreq <= '0';
      
    ELSIF clk80mhz'event AND clk80mhz = '1' THEN  -- rising clock edge
      s_wrreq_out   <= '0';
      rdreq_out     <= '0';
      busy          <= '0';                       -- default is "busy"
      trgFifo_rdreq <= '0';

      CASE TState IS

        -- wait for trigger
        WHEN SWaitTrig =>
          busy <= '1';                  -- "not busy" until trigger
          IF evt_trg = '1' THEN
            TState <= SFifoChk;
          END IF;

          -- only continue, if there is enough space in the upstream FIFO
        WHEN SFifoChk =>
          IF (NOT outfifo_almost_full) THEN
            TState <= STagWrd;
          END IF;

          -- strobe tag word into DDL Fifo
        WHEN STagWrd =>
          s_outdata   <= X"DEADFACE";
          s_wrreq_out <= '1';

          TState <= SRdSerA;

          -- deserialize the 16bit input stream into 32bit output
          -- words with appropriately timed write_request signals TO
          -- strobe the result into a FIFO.
          -- Stop when we see a word starting  with "0xE0" (the
          -- separator word generated by the 2nd cable on TCPU)
        WHEN SRdSerA =>
          rdreq_out <= '1';

          IF indata(15 DOWNTO 8) = X"E0" THEN
            block_end := true;
          END IF;

          IF fifo_empty = '0' THEN
            ctr                     := ctr + 1;
            s_outdata(15 DOWNTO 0)  <= indata;
            s_outdata(31 DOWNTO 16) <= s_outdata(15 DOWNTO 0);
          END IF;

          IF ctr = 2 THEN
            IF block_end THEN
              block_end := false;
              TState    <= SDelay;
            END IF;

            s_wrreq_out <= '1';
            ctr         := 0;
          END IF;

          delayCtr := 0;

          -- delay for a while (~13 us)
        WHEN SDelay =>
          delayCtr := delayCtr + 1;
          IF delayCtr = 1024 THEN
            TState <= SRdTrg;
          END IF;

          -- emtpy the trigger FIFO into the DDL FIFO 
        WHEN SRdTrg =>
          s_outdata(31 DOWNTO 20) <= X"A00";  -- trigger word
          s_outdata(19 DOWNTO 0)  <= trgFifo_q;

          trgFifo_rdreq <= '1';         -- NOT trgFifo_empty;
          s_wrreq_out   <= NOT trgFifo_empty;

          IF trgFifo_empty = '1' THEN
            TState <= SEnd;
          END IF;

          -- set up the "end" separator and strobe it into the FIFO
        WHEN SEnd =>
          s_outdata(31 DOWNTO 24) <= X"EA";
          s_outdata(23 DOWNTO 0)  <= (OTHERS => '0');
          s_wrreq_out             <= '1';

          TState <= SWaitTrig;          -- return to the beginning

        WHEN OTHERS =>
          TState <= SWaitTrig;
          
      END CASE;
      
    END IF;
  END PROCESS shifter;
  
END ARCHITECTURE a;
