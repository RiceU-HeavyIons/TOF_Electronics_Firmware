-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mux 

-- ============================================================
-- File Name: mux_2x32.vhd
-- Megafunction Name(s):
-- 			lpm_mux
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 4.1 Build 208 09/10/2004 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2004 Altera Corporation
--Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
--support information,  device programming or simulation file,  and any other
--associated  documentation or information  provided by  Altera  or a partner
--under  Altera's   Megafunction   Partnership   Program  may  be  used  only
--to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
--other  use  of such  megafunction  design,  netlist,  support  information,
--device programming or simulation file,  or any other  related documentation
--or information  is prohibited  for  any  other purpose,  including, but not
--limited to  modification,  reverse engineering,  de-compiling, or use  with
--any other  silicon devices,  unless such use is  explicitly  licensed under
--a separate agreement with  Altera  or a megafunction partner.  Title to the
--intellectual property,  including patents,  copyrights,  trademarks,  trade
--secrets,  or maskworks,  embodied in any such megafunction design, netlist,
--support  information,  device programming or simulation file,  or any other
--related documentation or information provided by  Altera  or a megafunction
--partner, remains with Altera, the megafunction partner, or their respective
--licensors. No other licenses, including any licenses needed under any third
--party's intellectual property, are provided herein.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY mux_2x32 IS
	PORT
	(
		data1x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data0x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		sel		: IN STD_LOGIC ;
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END mux_2x32;


ARCHITECTURE SYN OF mux_2x32 IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_2D (1 DOWNTO 0, 31 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT lpm_mux
	GENERIC (
		lpm_size		: NATURAL;
		lpm_widths		: NATURAL;
		lpm_width		: NATURAL;
		lpm_type		: STRING
	);
	PORT (
			sel	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			data	: IN STD_LOGIC_2D (1 DOWNTO 0, 31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	sub_wire5    <= data0x(31 DOWNTO 0);
	result    <= sub_wire0(31 DOWNTO 0);
	sub_wire1    <= sel;
	sub_wire2(0)    <= sub_wire1;
	sub_wire3    <= data1x(31 DOWNTO 0);
	sub_wire4(1, 0)    <= sub_wire3(0);
	sub_wire4(1, 1)    <= sub_wire3(1);
	sub_wire4(1, 2)    <= sub_wire3(2);
	sub_wire4(1, 3)    <= sub_wire3(3);
	sub_wire4(1, 4)    <= sub_wire3(4);
	sub_wire4(1, 5)    <= sub_wire3(5);
	sub_wire4(1, 6)    <= sub_wire3(6);
	sub_wire4(1, 7)    <= sub_wire3(7);
	sub_wire4(1, 8)    <= sub_wire3(8);
	sub_wire4(1, 9)    <= sub_wire3(9);
	sub_wire4(1, 10)    <= sub_wire3(10);
	sub_wire4(1, 11)    <= sub_wire3(11);
	sub_wire4(1, 12)    <= sub_wire3(12);
	sub_wire4(1, 13)    <= sub_wire3(13);
	sub_wire4(1, 14)    <= sub_wire3(14);
	sub_wire4(1, 15)    <= sub_wire3(15);
	sub_wire4(1, 16)    <= sub_wire3(16);
	sub_wire4(1, 17)    <= sub_wire3(17);
	sub_wire4(1, 18)    <= sub_wire3(18);
	sub_wire4(1, 19)    <= sub_wire3(19);
	sub_wire4(1, 20)    <= sub_wire3(20);
	sub_wire4(1, 21)    <= sub_wire3(21);
	sub_wire4(1, 22)    <= sub_wire3(22);
	sub_wire4(1, 23)    <= sub_wire3(23);
	sub_wire4(1, 24)    <= sub_wire3(24);
	sub_wire4(1, 25)    <= sub_wire3(25);
	sub_wire4(1, 26)    <= sub_wire3(26);
	sub_wire4(1, 27)    <= sub_wire3(27);
	sub_wire4(1, 28)    <= sub_wire3(28);
	sub_wire4(1, 29)    <= sub_wire3(29);
	sub_wire4(1, 30)    <= sub_wire3(30);
	sub_wire4(1, 31)    <= sub_wire3(31);
	sub_wire4(0, 0)    <= sub_wire5(0);
	sub_wire4(0, 1)    <= sub_wire5(1);
	sub_wire4(0, 2)    <= sub_wire5(2);
	sub_wire4(0, 3)    <= sub_wire5(3);
	sub_wire4(0, 4)    <= sub_wire5(4);
	sub_wire4(0, 5)    <= sub_wire5(5);
	sub_wire4(0, 6)    <= sub_wire5(6);
	sub_wire4(0, 7)    <= sub_wire5(7);
	sub_wire4(0, 8)    <= sub_wire5(8);
	sub_wire4(0, 9)    <= sub_wire5(9);
	sub_wire4(0, 10)    <= sub_wire5(10);
	sub_wire4(0, 11)    <= sub_wire5(11);
	sub_wire4(0, 12)    <= sub_wire5(12);
	sub_wire4(0, 13)    <= sub_wire5(13);
	sub_wire4(0, 14)    <= sub_wire5(14);
	sub_wire4(0, 15)    <= sub_wire5(15);
	sub_wire4(0, 16)    <= sub_wire5(16);
	sub_wire4(0, 17)    <= sub_wire5(17);
	sub_wire4(0, 18)    <= sub_wire5(18);
	sub_wire4(0, 19)    <= sub_wire5(19);
	sub_wire4(0, 20)    <= sub_wire5(20);
	sub_wire4(0, 21)    <= sub_wire5(21);
	sub_wire4(0, 22)    <= sub_wire5(22);
	sub_wire4(0, 23)    <= sub_wire5(23);
	sub_wire4(0, 24)    <= sub_wire5(24);
	sub_wire4(0, 25)    <= sub_wire5(25);
	sub_wire4(0, 26)    <= sub_wire5(26);
	sub_wire4(0, 27)    <= sub_wire5(27);
	sub_wire4(0, 28)    <= sub_wire5(28);
	sub_wire4(0, 29)    <= sub_wire5(29);
	sub_wire4(0, 30)    <= sub_wire5(30);
	sub_wire4(0, 31)    <= sub_wire5(31);

	lpm_mux_component : lpm_mux
	GENERIC MAP (
		lpm_size => 2,
		lpm_widths => 1,
		lpm_width => 32,
		lpm_type => "LPM_MUX"
	)
	PORT MAP (
		sel => sub_wire2,
		data => sub_wire4,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "2"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL result[31..0]
-- Retrieval info: USED_PORT: data1x 0 0 32 0 INPUT NODEFVAL data1x[31..0]
-- Retrieval info: USED_PORT: data0x 0 0 32 0 INPUT NODEFVAL data0x[31..0]
-- Retrieval info: USED_PORT: sel 0 0 0 0 INPUT NODEFVAL sel
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: CONNECT: @data 1 1 32 0 data1x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 0 32 0 data0x 0 0 32 0
-- Retrieval info: CONNECT: @sel 0 0 1 0 sel 0 0 0 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2x32.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2x32.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2x32.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2x32.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_2x32_inst.vhd TRUE
