mux_2to1_1bit_inst : mux_2to1_1bit PORT MAP (
		data1	 => data1_sig,
		data0	 => data0_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
