mux_2in_4bit_inst : mux_2in_4bit PORT MAP (
		data1x	 => data1x_sig,
		data0x	 => data0x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
