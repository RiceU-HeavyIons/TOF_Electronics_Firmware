SHIFTREG_inst : SHIFTREG PORT MAP (
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		shiftout	 => shiftout_sig
	);
